grammar lmlang;

nonterminal Type;

abstract production int_type
top::Type ::= 
{}

abstract production bool_type
top::Type ::= 
{}

abstract production module_type
top::Type ::=
{}

abstract production fun_type
top::Type ::=
{}

abstract production temp_type
top::Type ::=
{}