grammar scopegraphtest;
imports silver:testing;
mainTestSuite scopegraphtesting;