grammar scopetree;

global graphviz_font_size::String = "12";

function graphviz_draw_graph
String ::= graph::Graph<d r>
{
  return "";
}