grammar scope_tree_generic:ast;

{- Global label initialization -}

global mod_lab :: Label = mod_prod ();
global var_lab :: Label = var_prod ();
global rec_lab :: Label = rec_prod ();
global ext_lab :: Label = ext_prod ();
global imp_lab :: Label = imp_prod ();
global lex_lab :: Label = lex_prod ();

{- Global label order -}

global label_ord :: [[Label]] = [
  [mod_lab, var_lab, rec_lab],
  [ext_lab, imp_lab],
  [lex_lab]
];

{- Label equality -}

function label_eq
Boolean ::= l1::Label l2::Label
{
  return
    case (l1, l2) of
      (lex_prod (), lex_prod ()) -> true
    | (ext_prod (), ext_prod ()) -> true
    | (var_prod (), var_prod ()) -> true
    | (imp_prod (), imp_prod ()) -> true
    | (mod_prod (), mod_prod ()) -> true
    | (rec_prod (), rec_prod ()) -> true
    | _                            -> false
    end;
}

{- Labels -}

nonterminal Label;
synthesized attribute lab_str :: String occurs on Label;

abstract production lex_prod
top::Label ::= { top.lab_str = "LEX"; }

abstract production ext_prod
top::Label ::= { top.lab_str = "EXT"; }

abstract production var_prod
top::Label ::= { top.lab_str = "VAR"; }

abstract production imp_prod
top::Label ::= { top.lab_str = "IMP"; }

abstract production mod_prod
top::Label ::= { top.lab_str = "MOD"; }

abstract production rec_prod
top::Label ::= { top.lab_str = "REC"; }

{- Regular expressions -}

nonterminal Regex;
synthesized attribute nfa :: NFA occurs on Regex;

abstract production concatenate
top::Regex ::= r1::Regex r2::Regex
{ top.nfa = nfa_concatenate (r1.nfa, r2.nfa); }

abstract production star
top::Regex ::= r1::Regex
{ top.nfa = nfa_star (r1.nfa); }

abstract production alternate
top::Regex ::= r1::Regex r2::Regex
{ top.nfa = nfa_alternate (r1.nfa, r2.nfa); }

abstract production single
top::Regex ::= label::Label
{ top.nfa = nfa_single (label); }