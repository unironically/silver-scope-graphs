grammar scopegraph;