grammar scope_tree_generic:ast;

nonterminal Scope;