nonterminal LMR_Type;

abstract production rec_type
top::LMR_Type ::= s::Scope
{}