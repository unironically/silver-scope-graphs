grammar simple;

nonterminal Type;

abstract production int
top::Type ::=
{}

abstract production bool
top::Type ::=
{}

abstract production bottom
top::Type ::=
{}