grammar scopegraph;
