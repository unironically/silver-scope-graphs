grammar scopegraph;



------------------
-- Errors:
