grammar scope_tree_generic:ast;