grammar scopetree;