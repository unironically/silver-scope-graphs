grammar scopegraph_kw;